//=========================================================================
// Copyright (C) 2018 The C++ Component Model(COMO) Open Source Project
//
// Licensed under the Apache License, Version 2.0 (the "License");
// you may not use this file except in compliance with the License.
// You may obtain a copy of the License at
//
//      http://www.apache.org/licenses/LICENSE-2.0
//
// Unless required by applicable law or agreed to in writing, software
// distributed under the License is distributed on an "AS IS" BASIS,
// WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
// See the License for the specific language governing permissions and
// limitations under the License.
//=========================================================================

[
    uuid(42197c0a-0de1-4c11-8a35-4ed719e72695),
    uri("http://como.org/component/test/reflection/ReflectionTestUnit.so")
/*@
module ReflectionTestUnit FramacBlock ...
*/
]
module ReflectionTestUnit
{

include "ConstantTest.cdl"
include "MethodTest.cdl"

}
