//=========================================================================
// Copyright (C) 2021 The C++ Component Model(COMO) Open Source Project
//
// Licensed under the Apache License, Version 2.0 (the "License");
// you may not use this file except in compliance with the License.
// You may obtain a copy of the License at
//
//      http://www.apache.org/licenses/LICENSE-2.0
//
// Unless required by applicable law or agreed to in writing, software
// distributed under the License is distributed on an "AS IS" BASIS,
// WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
// See the License for the specific language governing permissions and
// limitations under the License.
//=========================================================================


namespace como {

[
    uuid(00000000-0000-0000-0000-000000000101),
    version(0.1.0)
]
interface IComoFunctionSafetyObject
{
    const Integer CFSO_ExpireVALID = 0;
    const Integer CFSO_ExpireTime = 1;

    IsValid(
        [out] Integer& isValid);

    InvalidObject(
        [in] Integer isValid);

    GetChecksum(
        [out] Long& lastChecksum,
        [out] Long& currentChecksum);
}

}
