//=========================================================================
// Copyright (C) 2018 The C++ Component Model(COMO) Open Source Project
//
// Licensed under the Apache License, Version 2.0 (the "License");
// you may not use this file except in compliance with the License.
// You may obtain a copy of the License at
//
//      http://www.apache.org/licenses/LICENSE-2.0
//
// Unless required by applicable law or agreed to in writing, software
// distributed under the License is distributed on an "AS IS" BASIS,
// WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
// See the License for the specific language governing permissions and
// limitations under the License.
//=========================================================================

include "ICelestialBody.cdl"

interface Universe::IPlanet;

namespace Universe {

[
    uuid(c2d17b6c-8dd8-42cb-8aae-6f035ae9ecc8),
    version(0.1.0)
]
interface ISatellite : ICelestialBody
{
    const CelestialBodyKind KIND = satellite;

    GetAroundPlanet(
        [out] IPlanet** planet);

    GetDistanceToPlanet(
        [out] Double* distance);

    GetOrbitalPeriod(
        [out] Integer* hours);
}

} // namespace Universe
