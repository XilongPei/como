//=========================================================================
// Copyright (C) 2018 The C++ Component Model(COMO) Open Source Project
//
// Licensed under the Apache License, Version 2.0 (the "License");
// you may not use this file except in compliance with the License.
// You may obtain a copy of the License at
//
//      http://www.apache.org/licenses/LICENSE-2.0
//
// Unless required by applicable law or agreed to in writing, software
// distributed under the License is distributed on an "AS IS" BASIS,
// WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
// See the License for the specific language governing permissions and
// limitations under the License.
//=========================================================================

interface como::io::ISerializable;

namespace como {
namespace core {

[
    uuid(df471c09-381f-40c4-9e24-c92b31dd9146),
    version(0.1.0)
]
coclass CBoolean
{
    Constructor(
           [in] Boolean value);

   interface IBoolean;
   interface ISerializable;
   interface IComparable;
}

[
    uuid(bdf665c0-8a7a-4621-ba55-e6a097dfc85d),
    version(0.1.0)
]
coclass CByte
{
    Constructor(
        [in] Byte value);

    interface IByte;
    interface INumber;
    interface ISerializable;
    interface IComparable;
}

[
    uuid(f30fd610-ee65-4fc0-8191-e840c7f73125),
    version(0.1.0)
]
coclass CChar
{
    Constructor(
        [in] Char value);

    interface IChar;
    interface ISerializable;
    interface IComparable;
}

[
    uuid(38abe6d2-1428-4a97-8177-b24d09593d15),
    version(0.1.0)
]
coclass CDouble
{
    Constructor(
        [in] Double value);

    interface IDouble;
    interface INumber;
    interface ISerializable;
    interface IComparable;
}

[
    uuid(569b10e8-38d5-41f6-a89a-36fcde449413),
    version(0.1.0)
]
coclass CFloat
{
    Constructor(
        [in] Float value);

    interface IFloat;
    interface INumber;
    interface ISerializable;
    interface IComparable;
}

[
    uuid(55469170-d13e-4567-9435-3bf4c5ebf1e4),
    version(0.1.0)
]
coclass CInteger
{
    Constructor(
        [in] Integer value);

    interface IInteger;
    interface INumber;
    interface ISerializable;
    interface IComparable;
}

[
    uuid(bc8830e2-23f7-4a25-b61e-dbc9cce385b2),
    version(0.1.0)
]
coclass CLong
{
    Constructor(
        [in] Long value);

    interface ILong;
    interface INumber;
    interface ISerializable;
    interface IComparable;
}

[
    uuid(cdff023b-ba1b-4e14-bf1b-8ebf9fe80214),
    version(0.1.0)
]
coclass CShort
{
    Constructor(
        [in] Short value);

    interface IShort;
    interface INumber;
    interface ISerializable;
    interface IComparable;
}

[
    uuid(16a75841-ffee-43a5-bd5c-4f8362361b35),
    version(0.1.0)
]
coclass CStackTrace
{
    Constructor();

    Constructor(
        [in] String message);

    interface IStackTrace;
    interface ISerializable;
}

[
    uuid(c2fee305-a2bb-453a-9248-473bbef55fd0),
    version(0.1.0)
]
coclass CStackTraceElement
{
    Constructor(
        [in] Integer no,
        [in] HANDLE  pc,
        [in] String  soname,
        [in] String  symbol,
        [in] HANDLE  relOffset,
        [in] HANDLE  thisPointer);

    interface IStackTraceElement;
    interface ISerializable;
}

[
    uuid(10e6419e-b8d0-44be-b309-54086eb3e560),
    version(0.1.0)
]
coclass CString
{
    Constructor(
        [in] String str);

    interface ISerializable;
    interface ICharSequence;
    interface IComparable;
    interface IString;
}

[
    uuid(8c3a55f1-63c5-4abd-b68c-46773877a655),
    version(0.1.0)
]
coclass CStringBuffer
{
    Constructor();

    Constructor(
        [in] Integer capacity);

    Constructor(
        [in] String str);

    Constructor(
        [in] ICharSequence* seq);

    interface ISerializable;
    interface ICharSequence;
    interface IStringBuffer;
}

[
    uuid(cbc6b55a-c06e-4ddc-b7f8-f0cc0bf94ff9),
    version(0.1.0)
]
coclass CStringBuilder
{
    Constructor();

    Constructor(
        [in] Integer capacity);

    Constructor(
        [in] String str);

    Constructor(
        [in] ICharSequence* seq);

    interface ISerializable;
    interface ICharSequence;
    interface IStringBuilder;
}

}
}
