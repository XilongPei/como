//=========================================================================
// Copyright (C) 2018 The C++ Component Model(COMO) Open Source Project
//
// Licensed under the Apache License, Version 2.0 (the "License");
// you may not use this file except in compliance with the License.
// You may obtain a copy of the License at
//
//      http://www.apache.org/licenses/LICENSE-2.0
//
// Unless required by applicable law or agreed to in writing, software
// distributed under the License is distributed on an "AS IS" BASIS,
// WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
// See the License for the specific language governing permissions and
// limitations under the License.
//=========================================================================

namespace como {
namespace test {
namespace rpc {

enum TestEnum 
{
    Monday,
    Tuesday,
    Wednesday,
    Thursday,
    Friday,
    Saturday,
    Sunday
}

[
    uuid(ae56a8d1-28a5-eca7-a578-97ebbf8bba6e),
    version(0.1.0)
]
interface IService2
{
    TestMethod1(
        [in] Array<Integer> arg1,
        [out] Array<Integer>* result1);

    TestMethod2(
        [in] Integer arg1,
        [out] Char* result1,
        [out] Char* result2,
        [out] Char* result3,
        [out] Char* result4);

    TestMethod3(
        [in] TestEnum arg1,
        [out] String& result1);

    TestMethod4(
        [in] Triple arg1,
        [out] Char* result1,
        [out] Long& result2,
        [out] TypeKind& result3);
}

[
    uuid(181919c5-e8b6-ef7a-31e5-a298e0f1eb9c),
    version(0.1.0)
]
coclass CService2
{
    interface IService2;
}

}
}
}