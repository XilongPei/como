//=========================================================================
// Copyright (C) 2024 The C++ Component Model(COMO) Open Source Project
//
// Licensed under the Apache License, Version 2.0 (the "License");
// you may not use this file except in compliance with the License.
// You may obtain a copy of the License at
//
//      http://www.apache.org/licenses/LICENSE-2.0
//
// Unless required by applicable law or agreed to in writing, software
// distributed under the License is distributed on an "AS IS" BASIS,
// WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
// See the License for the specific language governing permissions and
// limitations under the License.
//=========================================================================

namespace como {
namespace test {
namespace reflection {

[
    uuid(6611bd57-14c2-4b5f-b971-9d47b122fc22),
    version(0.1.0)
]
interface IMethodTest2
{
    TestMethod1(
        [in] Integer arg,
        [out] Integer& result);

    TestMethod2(
        [in] Float arg,
        [out] Float& result);
}

[
    uuid(85511188-d0e5-42b0-99d7-483a0129ac95),
    version(0.1.0),
    FuncSafetySetting("expire")
]
coclass CMethodTester2
{
    interface IMethodTest2;
    interface IObjectObserver;
}

}
}
}
