//=========================================================================
// Copyright (C) 2018 The C++ Component Model(COMO) Open Source Project
//
// Licensed under the Apache License, Version 2.0 (the "License");
// you may not use this file except in compliance with the License.
// You may obtain a copy of the License at
//
//      http://www.apache.org/licenses/LICENSE-2.0
//
// Unless required by applicable law or agreed to in writing, software
// distributed under the License is distributed on an "AS IS" BASIS,
// WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
// See the License for the specific language governing permissions and
// limitations under the License.
//=========================================================================

namespace como {

enum RPCType
{
    Local,
    Remote
}

enum RPCPeer
{
    Proxy,
    Stub
}

[
    uuid(3d29cb55-f7d1-4b79-9e63-ad14a57fd9f1),
    version(0.1.0)
]
interface IParcel
{
    ReadChar(
        [out] Char& value);

    WriteChar(
        [in] Char value);

    ReadByte(
        [out] Byte& value);

    WriteByte(
        [in] Byte value);

    ReadShort(
        [out] Short& value);

    WriteShort(
        [in] Short value);

    ReadInteger(
        [out] Integer& value);

    WriteInteger(
        [in] Integer value);

    ReadLong(
        [out] Long& value);

    WriteLong(
        [in] Long value);

    ReadFloat(
        [out] Float& value);

    WriteFloat(
        [in] Float value);

    ReadDouble(
        [out] Double& value);

    WriteDouble(
        [in] Double value);

    ReadBoolean(
        [out] Boolean& value);

    WriteBoolean(
        [in] Boolean value);

    ReadString(
        [out] String& value);

    WriteString(
        [in] String value);

    ReadCoclassID(
        [out] CoclassID& value);

    WriteCoclassID(
        [in] CoclassID value);

    ReadComponentID(
        [out] ComponentID& value);

    WriteComponentID(
        [in] ComponentID value);

    ReadInterfaceID(
        [out] InterfaceID& value);

    WriteInterfaceID(
        [in] InterfaceID value);

    ReadECode(
        [out] ECode& value);

    WriteECode(
        [in] ECode value);

    ReadEnumeration(
        [out] Integer& value);

    WriteEnumeration(
        [in] Integer value);

    ReadArray(
        [out] Triple* array);

    WriteArray(
        [in] Triple array);

    ReadInterface(
        [out] IInterface&& value);

    WriteInterface(
        [in] IInterface* value);

    GetData(
        [out] HANDLE& data);

    GetDataSize(
        [out] Long& size);

    SetData(
        [in] HANDLE data,
        [in] Long size);

    GetDataPosition(
        [out] Long& pos);

    SetDataPosition(
        [in] Long pos);

    GetPayload(
        [out] HANDLE& payload);

    SetPayload(
        [in] HANDLE payload,
        [in] Boolean release);
}

[
    uuid(6abf4491-874b-4e8c-855b-d74f2e20cf6b),
    version(0.1.0)
]
interface IParcelable
{
    ReadFromParcel(
        [in] IParcel* source);

    WriteToParcel(
        [in] IParcel* dest);
}

[
    uuid(84ee26c6-6c0a-4329-b627-54e5fc3b06a8),
    version(0.1.0)
]
interface IInterfacePack
{
    GetCoclassID(
        [out] CoclassID& cid);

    GetInterfaceID(
        [out] InterfaceID& iid);

    IsParcelable(
        [out] Boolean& parcelable);

    SetServerName(
        [in] String serverName);

    GetServerName(
        [out] String& serverName);

    GetHashCode(
        [out] Integer& hash);

    GetServerIdString(
        [out] String& serverIdString);
}

interface IArgumentList;
interface IDeathRecipient;
interface IMetaMethod;
interface IProxy;
interface IStub;

[
    uuid(bf89f2ce-ba5f-4f5d-a866-9e34048ee009),
    version(0.1.0)
]
interface IRPCChannel
{
    Apply(
        [in] IInterfacePack* ipack);

    GetRPCType(
        [out] RPCType& type);

    GetServerName(
        [out] String& serverName);

    SetServerName(
        [in] String serverName);

    IsPeerAlive(
        [out] Boolean& alive);

    ReleasePeer(
        [out] Boolean& alive);

    LinkToDeath(
        [in] IProxy* proxy,
        [in] IDeathRecipient* recipient,
        [in] HANDLE cookie = 0,
        [in] Integer flags = 0);

    UnlinkToDeath(
        [in] IProxy* proxy,
        [in] IDeathRecipient* recipient,
        [in] HANDLE cookie = 0,
        [in] Integer flags = 0,
        [out] IDeathRecipient&* outRecipient = nullptr);

    GetComponentMetadata(
        [in] CoclassID cid,
        [out, callee] Array<Byte>& metadata);

    Invoke(
        [in] IMetaMethod* method,
        [in] IParcel* argParcel,
        [out] IParcel&& resParcel);

    StartListening(
        [in] IStub* stub);

    Match(
        [in] IInterfacePack* ipack,
        [out] Boolean& matched);
}

[
    uuid(d1adf1f9-2062-45fd-aa33-edd481a04417),
    version(0.1.0)
]
interface IRPCChannelFactory
{
    CreateInterfacePack(
        [out] IInterfacePack&& ipack);

    CreateParcel(
        [out] IParcel&& parcel);

    CreateChannel(
        [in] RPCPeer peer,
        [out] IRPCChannel&& channel);

    MarshalInterface(
        [in] IInterface* object,
        [out] IInterfacePack&& ipack);

    UnmarshalInterface(
        [in] IInterfacePack* data,
        [out] IInterface&& object);
}

[
    uuid(2598f97d-0e6b-45a2-8c21-ffeca8347233),
    version(0.1.0)
]
interface IProxy
{
    GetTargetCoclass(
        [out] IMetaCoclass&& target);

    IsStubAlive(
        [out] Boolean& alive);

    ReleaseStub(
        [out] Boolean& alive);

    LinkToDeath(
        [in] IDeathRecipient* recipient,
        [in] HANDLE cookie = 0,
        [in] Integer flags = 0);

    UnlinkToDeath(
        [in] IDeathRecipient* recipient,
        [in] HANDLE cookie = 0,
        [in] Integer flags = 0,
        [out] IDeathRecipient&* outRecipient = nullptr);
}

[
    uuid(2598f97d-0e6b-45a2-8c21-ffeca8347233),
    version(0.1.0)
]
interface IDeathRecipient
{
    StubDied(
        [in] IProxy* who);
}

[
    uuid(7752e566-880a-4abd-99b9-417176e0644f),
    version(0.1.0)
]
interface IStub
{
    Match(
        [in] IInterfacePack* ipack,
        [out] Boolean& matched);

    Invoke(
        [in] IParcel* argParcel,
        [out] IParcel&& resParcel);
}

}
