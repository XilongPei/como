//=========================================================================
// Copyright (C) 2024 The C++ Component Model(COMO) Open Source Project
//
// Licensed under the Apache License, Version 2.0 (the "License");
// you may not use this file except in compliance with the License.
// You may obtain a copy of the License at
//
//      http://www.apache.org/licenses/LICENSE-2.0
//
// Unless required by applicable law or agreed to in writing, software
// distributed under the License is distributed on an "AS IS" BASIS,
// WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
// See the License for the specific language governing permissions and
// limitations under the License.
//=========================================================================

namespace como {
namespace test {
namespace reflection {

[
    uuid(6611bd57-14c2-4b5f-b971-9d47b122fc21),
    version(0.1.0)
/*@
$$$ interface IMethodTest FramacBlock ... $$$
*/
]
interface IMethodTest
{
    TestMethod1(
        [in] Integer arg,
        [out] Integer& result);

/*@
$$$ TestMethod2 FramacBlock ... $$$
*/
    TestMethod2(
        [in] Float arg,
        [out] Float& result);

    TestMethod3(
        [in] Integer arg1,
        [in] Long arg2,
        [in] Boolean arg3,
        [in] Char arg4,
        [in] Short arg5,
        [in] Integer arg6);

    TestMethod4(
        [in] Integer arg1,
        [in] Long arg2,
        [in] Boolean arg3,
        [in] Char arg4,
        [in] Short arg5,
        [in] Double arg6,
        [in] Float arg7,
        [in] Integer arg8,
        [out] Double& result);

    TestMethod5(
        [in] Integer arg1,
        [in] Long arg2,
        [in] Boolean arg3,
        [in] Char arg4,
        [in] Short arg5,
        [in] Double arg6,
        [in] Float arg7,
        [in] Integer arg8,
        [in] Float arg9,
        [in] Double arg10,
        [in] Double arg11,
        [in] Float arg12,
        [in] Float arg13,
        [in] Double arg14,
        [in] Double arg15,
        [in] Float arg16,
        [out] Double& result);

    TestMethod6(
        [in] Integer arg1,
        [in] Long arg2,
        [in] Boolean arg3,
        [in] Char arg4,
        [in] Short arg5,
        [in] Double arg6,
        [in] Float arg7,
        [in] Integer arg8,
        [in] Float arg9,
        [in] Double arg10,
        [in] Double arg11,
        [in] Float arg12,
        [in] Float arg13,
        [in] Double arg14,
        [in] Double arg15,
        [in] Float arg16,
        [out] Integer& result1,
        [out] Double& result2);
}

[
    uuid(85511188-d0e5-42b0-99d7-483a0129ac94),
    version(0.1.0),
    FuncSafetySetting("expire")
]
coclass CMethodTester
{
    //interface IComoFunctionSafetyObject;
    interface IMethodTest;
    interface IObjectObserver;
}

}
}
}
