//=========================================================================
// Copyright (C) 2018 The C++ Component Model(COMO) Open Source Project
//
// Licensed under the Apache License, Version 2.0 (the "License");
// you may not use this file except in compliance with the License.
// You may obtain a copy of the License at
//
//      http://www.apache.org/licenses/LICENSE-2.0
//
// Unless required by applicable law or agreed to in writing, software
// distributed under the License is distributed on an "AS IS" BASIS,
// WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
// See the License for the specific language governing permissions and
// limitations under the License.
//=========================================================================

include "ISolarSystemPlanet.cdl"
include "IMoon.cdl"

namespace Universe {
namespace MilkyWay {
namespace SolarSystem {

[
    uuid(53b51043-e26f-44d6-84cf-094a5fade941),
    version(0.1.0)
]
interface IEarth : ISolarSystemPlanet
{
    const Double WEIGHT = 5.972e24;

    GetDistanceToMoon(
        [out] Double* distance);
}

} // namespace SolarSystem
} // namespace MilkyWay
} // namespace Universe
