//=========================================================================
// Copyright (C) 2018 The C++ Component Model(COMO) Open Source Project
//
// Licensed under the Apache License, Version 2.0 (the "License");
// you may not use this file except in compliance with the License.
// You may obtain a copy of the License at
//
//      http://www.apache.org/licenses/LICENSE-2.0
//
// Unless required by applicable law or agreed to in writing, software
// distributed under the License is distributed on an "AS IS" BASIS,
// WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
// See the License for the specific language governing permissions and
// limitations under the License.
//=========================================================================

/**
 * ISolarSystemPlanet is an IPlanet in solar system.
 */

include "IPlanet.cdl"

namespace Universe {
namespace MilkyWay {
namespace SolarSystem {

[
    uuid(768600c6-0f61-40ca-80a3-ccdc0c09c54e),
    version(0.1.0),
    description("This is the definiton of ISolarSystemPlanet.")
]
interface ISolarSystemPlanet : IPlanet
{
    const String STAR_NAME = "Sun";

    GetDistanceToSun(
        [out] Double* distance);
}

} // namespace SolarSystem
} // namespace MilkyWay
} // namespace Universe
